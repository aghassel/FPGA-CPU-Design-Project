module alu #(parameter wordSize = 32)(
    input clk, clr, read, MDRin,
    input [wordSize-1:0] BusMuxOut, Mdatain,
    output reg [31:0] Q
);

endmodule