`timescale 1ns/1ps

module ctrl_unit;



end module 