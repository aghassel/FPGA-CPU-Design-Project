//refer to diagram, get inputs for R0signal and for the contents of R0 (acc registers)
module bus  #(parameter wordSize = 32)(
    input R0out, R1out, R2out, R3out, R4out, R5out, R6out, R7out, R8out, R9out, R10out, R11out, R12out, R13out, R14out, R15out,
    input HIout, LOout, Zhighout, Zlowout, PCout, MDRout, InPortout, Cout,
    input [wordSize-1:0] BusMuxIn_R0, BusMuxIn_R1, BusMuxIn_BusMuxIn_R2, BusMuxIn_R3, BusMuxIn_R4, BusMuxIn_R5, BusMuxIn_R6, BusMuxIn_R7, BusMuxIn_R8, BusMuxIn_R9, BusMuxIn_R10, BusMuxIn_R11, BusMuxIn_R12, BusMuxIn_R13, BusMuxIn_R14, BusMuxIn_R15,
    input [wordSize-1:0] BusMuxIn_HI, BusMuxIn_LO, BusMuxIn_Zhigh, BusMuxIn_Zlow, BusMuxIn_PC, BusMuxIn_MDR, BusMuxIn_InPort
    output reg [wordSize-1:0] BusMuxOut
);

wire [5:0] s;

wire [wordSize-1:0] c_sign_extended;

assign c_sign_extended = (Cout == 0) ? 32'd0 : 32'd1;

encoder32to5 myEncoder(
//input wire [31:0]ein, output reg [4:0] eout
.ein[0](R0out),
.ein[1](R1out),
.ein[2](R2out),
.ein[3](R3out),
.ein[4](R4out),
.ein[5](R5out),
.ein[6](R6out),
.ein[7](R7out),
.ein[8](R8out),
.ein[9](R9out),
.ein[10](R10out),
.ein[11](R11out),
.ein[12](R12out),
.ein[13](R13out),
.ein[14](R14out),
.ein[15](R15out),
.ein[16](HIout),
.ein[17](LOout),
.ein[18](Zhighout),
.ein[19](Zlowout),
.ein[20](PCout),
.ein[21](MDRout),
.ein[22](InPortout),
.ein[23](Cout),
.ein[24](0),
.ein[25](0),
.ein[26](0),
.ein[27](0),
.ein[28](0),
.ein[29](0),
.ein[30](0),
.ein[31](0),
.eout(s)
);

mux32to1 BusMux(
    /*
    input wire [31:0] data0, data1, data2, data3, data4, data5, data6, data7, data8, data9, data10, data11, data12, data13, data14, data15, data16, data17, data18, data19, data20, data21, data22, data23, data24, data25, data26, data27, data28, data29, data30, data31;
	input wire [4:0] s;
	output reg [31:0] out;
    */
    .data0(BusMuxIn_R0),
    .data1(BusMuxIn_R1),
    .data2(BusMuxIn_R2),
    .data3(BusMuxIn_R3),
    .data4(BusMuxIn_R4),
    .data5(BusMuxIn_R5),
    .data6(BusMuxIn_R6),
    .data7(BusMuxIn_R7),
    .data8(BusMuxIn_R8),
    .data9(BusMuxIn_R9),
    .data10(BusMuxIn_R10),
    .data11(BusMuxIn_R11),
    .data12(BusMuxIn_R12),
    .data13(BusMuxIn_R13),
    .data14(BusMuxIn_R14),
    .data15(BusMuxIn_R15),
    .data16(BusMuxIn_HI),
    .data17(BusMuxIn_LO),
    .data18(BusMuxIn_Zhigh),
    .data19(BusMuxIn_Zlow),
    .data20(BusMuxIn_PC),
    .data21(BusMuxIn_MDR),
    .data22(BusMuxIn_InPort),
    .data23(c_sign_extended),
    .data24(0),
    .data25(0),
    .data26(0),
    .data27(0),
    .data28(0),
    .data29(0),
    .data30(0),
    .data31(0),
    .s(s),
    .out(BusMuxOut)
    );
    
    endmodule