//bussy module

module bus  #(parameter wordSize = 32)(
    input wire [14:0] r_x,
    input regLOout,
    input Zhighout,
    input Zlowout,
    input PCout,
    input 
//incomplete - reworking components
)

endmodule